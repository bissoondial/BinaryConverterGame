module lightblinker (input clk, input [7:0] number, output [7:0] lights);

assign lights = number;

endmodule